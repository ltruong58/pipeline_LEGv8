//////////////////////////////////////////////////////////////////////////////////
//										
// 64-bit Mux							
// 										
//////////////////////////////////////////////////////////////////////////////////

module FullMux(
	input [63:0] a, b,
	input select,
	output [63:0] out
	);

	assign out = (select == 0) ?  a : b;

endmodule